module DCS(
    input a,
    input b,
    output f,
    output f1
);
assign f = a^b;
assign f1 = 1'b1;
endmodule
